// Level 3: Deepest level - simple value macros
`define LEVEL3_MACRO 3
`define DEEP_MACRO 42
