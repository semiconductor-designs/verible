// Test case for STR_003: Deep hierarchy (>5 levels of instantiation)
// Note: Full test would require actual deep nesting

module str_deep_hierarchy_violation;
  // STR_003: Simulated deep hierarchy marker
  // Real implementation would analyze actual instantiation depth
  // For testing, we use a comment marker
  // hierarchy:depth=6
  
  logic clk, data;
endmodule

