// Empty module with no ports

module empty_module;
  // No ports
endmodule

module top;
  empty_module u_empty();
endmodule

