// Test case: Empty module with no functions
module empty_module (
  input logic clk
);
  // No functions or tasks defined
endmodule

