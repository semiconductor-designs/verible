// Level 1: Includes level 2
`include "level2.svh"

// Additional macro at this level
`define LEVEL1_MACRO 1
