// Level 2: Includes level 3
`include "level3.svh"

// Additional macro at this level
`define LEVEL2_MACRO 2
