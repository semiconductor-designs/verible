// Copyright 2025 The Verible Authors.
// Edge case: Minimal 1-line module (buffer)
module str_edge_minimal_1line (input wire d, output wire q); assign q = d; endmodule

