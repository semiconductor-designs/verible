// Empty module (edge case)
module empty_module (
  input  logic clk
);
  
  // No signals, no data flow
  // This tests handling of empty modules
  
endmodule

