// Test case for NAM_001: Module naming convention
// Convention: module names should be lowercase with underscores (snake_case)

// Violation: PascalCase
module MyModule;
endmodule

// Violation: camelCase
module myFancyModule;
endmodule

// Good: snake_case
module my_good_module;
endmodule

